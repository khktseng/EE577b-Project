module mac_units(
	input clk,
	input reset,

