module divider(
	input [0:63] op1, op2,
	input [1:0] ww,
	output [0:63] mul_out
	);

endmodule
