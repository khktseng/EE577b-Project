// cardinal NOC verilog

module gold_router(
	input clk, reset,
	output polarity,

	input cwsi, ccwsi, pesi,
	output cwri, ccwri, peri,
	input [63:0] cwdi, ccwdi, pedi,

	output cwso, ccwso, peso,
	input cwro, ccwro, pero,
	output [63:0] cwdo, ccwdo, pedo
	);

	



endmodule
